module tb_simulation;
// signals to be connected between image_read and image_write modules
reg HCLK, HRESETn;
wire          data_write;
wire [ 7 : 0] data_R0;
wire [ 7 : 0] data_G0;
wire [ 7 : 0] data_B0;
wire [ 7 : 0] data_R1;
wire [ 7 : 0] data_G1;
wire [ 7 : 0] data_B1;
wire enc_done;
wire write_done;
//--------------------------------------------------------------------------------------------------------------
//start your code here...

endmodule
